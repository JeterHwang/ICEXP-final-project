module ALUlev1_tb;
    input [63:0] 
endmodule