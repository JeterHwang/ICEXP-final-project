module ALU_tb;
    reg clk;
    reg rst_n;
    reg [31:0] mat_in;
    reg [31:0] vec_in;
    reg [3:0] ipv_in;

     
endmodule